module tdc_top (
    
);

endmodule //tdc_top