library verilog;
use verilog.vl_types.all;
entity tb_spad is
end tb_spad;
