module decode (
    input  wire [31:0]  data_in,
    output reg  [ 4:0]  data_out
);

always @(*) begin
    case (data_in)
    0_1111_1111_1111_111:    data_out = 5'b0_0000; 
    0_0111_1111_1111_111:    data_out = 5'b0_0001; 
    0_0011_1111_1111_111:    data_out = 5'b0_0010; 
    0_0001_1111_1111_111:    data_out = 5'b0_0011; 
    0_0000_1111_1111_111:    data_out = 5'b0_0100; 
    0_0000_0111_1111_111:    data_out = 5'b0_0101; 
    0_0000_0011_1111_111:    data_out = 5'b0_0110; 
    0_0000_0001_1111_111:    data_out = 5'b0_0111; 

    0_0000_0000_1111_111:    data_out = 5'b0_1000; 
    0_0000_0000_0111_111:    data_out = 5'b0_1001; 
    0_0000_0000_0011_111:    data_out = 5'b0_1010; 
    0_0000_0000_0001_111:    data_out = 5'b0_1011; 
    0_0000_0000_0000_111:    data_out = 5'b0_1100; 
    0_0000_0000_0000_011:    data_out = 5'b0_1101; 
    0_0000_0000_0000_001:    data_out = 5'b0_1110; 
    0_0000_0000_0000_000:    data_out = 5'b0_1111; 

    1_0000_0000_0000_000:    data_out = 5'b1_0000;   
    1_1000_0000_0000_000:    data_out = 5'b1_0001; 
    1_1100_0000_0000_000:    data_out = 5'b1_0010; 
    1_1110_0000_0000_000:    data_out = 5'b1_0011; 
    1_1111_0000_0000_000:    data_out = 5'b1_0100; 
    1_1111_1000_0000_000:    data_out = 5'b1_0101; 
    1_1111_1100_0000_000:    data_out = 5'b1_0110; 
    1_1111_1110_0000_000:    data_out = 5'b1_0111; 

    1_1111_1111_0000_000:    data_out = 5'b1_1000; 
    1_1111_1111_1000_000:    data_out = 5'b1_1001; 
    1_1111_1111_1100_000:    data_out = 5'b1_1010; 
    1_1111_1111_1110_000:    data_out = 5'b1_1011; 
    1_1111_1111_1111_000:    data_out = 5'b1_1100; 
    1_1111_1111_1111_100:    data_out = 5'b1_1101; 
    1_1111_1111_1111_110:    data_out = 5'b1_1110; 
    1_1111_1111_1111_111:    data_out = 5'b1_1111; 

    default: data_out = 5'b0_0000;
    endcase
end
    0100 0000 0000 0000:    data_out = 5'b0_0000; 
    0010 0000 0000 0000:    data_out = 5'b0_0001; 
    0001 0000 0000 0000:    data_out = 5'b0_0010; 
    0000 1000 0000 0000:    data_out = 5'b0_0011; 
    0000 0100 0000 0000:    data_out = 5'b0_0100; 
    0000 0010 0000 0000:    data_out = 5'b0_0101; 
    0000 0001 0000 0000:    data_out = 5'b0_0110; 
    0000 0000 1000 0000:    data_out = 5'b0_0111; 

    0000 0000 0100 0000:    data_out = 5'b0_1000; 
    0000 0000 0010 0000:    data_out = 5'b0_1001; 
    0000 0000 0001 0000:    data_out = 5'b0_1010; 
    0000 0000 0000 1000:    data_out = 5'b0_1011; 
    0000 0000 0000 0100:    data_out = 5'b0_1100; 
    0000 0000 0000 0010:    data_out = 5'b0_1101; 
    0000 0000 0000 0001:    data_out = 5'b0_1110; 
    1000 0000 0000 0000:    data_out = 5'b0_1111;  

endmodule //decode