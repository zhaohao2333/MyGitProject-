module decode (
    input  wire [31:0]  data_in,
    output reg  [ 4:0]  data_out
);

always @(*) begin
    case (data_in)
    32'b0000_0000_0000_0000_1111_1111_1111_1111:    data_out = 5'b0_0000; 
    32'b1000_0000_0000_0000_0111_1111_1111_1111:    data_out = 5'b0_0001; 
    32'b1100_0000_0000_0000_0011_1111_1111_1111:    data_out = 5'b0_0010; 
    32'b1110_0000_0000_0000_0001_1111_1111_1111:    data_out = 5'b0_0011; 
    32'b1111_0000_0000_0000_0000_1111_1111_1111:    data_out = 5'b0_0100; 
    32'b1111_1000_0000_0000_0000_0111_1111_1111:    data_out = 5'b0_0101; 
    32'b1111_1100_0000_0000_0000_0011_1111_1111:    data_out = 5'b0_0110; 
    32'b1111_1110_0000_0000_0000_0001_1111_1111:    data_out = 5'b0_0111; 

    32'b1111_1111_0000_0000_0000_0000_1111_1111:    data_out = 5'b0_1000; 
    32'b1111_1111_1000_0000_0000_0000_0111_1111:    data_out = 5'b0_1001; 
    32'b1111_1111_1100_0000_0000_0000_0011_1111:    data_out = 5'b0_1010; 
    32'b1111_1111_1110_0000_0000_0000_0001_1111:    data_out = 5'b0_1011; 
    32'b1111_1111_1111_0000_0000_0000_0000_1111:    data_out = 5'b0_1100; 
    32'b1111_1111_1111_1000_0000_0000_0000_0111:    data_out = 5'b0_1101; 
    32'b1111_1111_1111_1100_0000_0000_0000_0011:    data_out = 5'b0_1110; 
    32'b1111_1111_1111_1110_0000_0000_0000_0001:    data_out = 5'b0_1111;
    
    32'b1111_1111_1111_1111_0000_0000_0000_0000:    data_out = 5'b1_0000;   
    32'b0111_1111_1111_1111_1000_0000_0000_0000:    data_out = 5'b1_0001; 
    32'b0011_1111_1111_1111_1100_0000_0000_0000:    data_out = 5'b1_0010; 
    32'b0001_1111_1111_1111_1110_0000_0000_0000:    data_out = 5'b1_0011; 
    32'b0000_1111_1111_1111_1111_0000_0000_0000:    data_out = 5'b1_0100; 
    32'b0000_0111_1111_1111_1111_1000_0000_0000:    data_out = 5'b1_0101; 
    32'b0000_0011_1111_1111_1111_1100_0000_0000:    data_out = 5'b1_0110; 
    32'b0000_0001_1111_1111_1111_1110_0000_0000:    data_out = 5'b1_0111; 

    32'b0000_0000_1111_1111_1111_1111_0000_0000:    data_out = 5'b1_1000; 
    32'b0000_0000_0111_1111_1111_1111_1000_0000:    data_out = 5'b1_1001; 
    32'b0000_0000_0011_1111_1111_1111_1100_0000:    data_out = 5'b1_1010; 
    32'b0000_0000_0001_1111_1111_1111_1110_0000:    data_out = 5'b1_1011; 
    32'b0000_0000_0000_1111_1111_1111_1111_0000:    data_out = 5'b1_1100; 
    32'b0000_0000_0000_0111_1111_1111_1111_1000:    data_out = 5'b1_1101; 
    32'b0000_0000_0000_0011_1111_1111_1111_1100:    data_out = 5'b1_1110; 
    32'b0000_0000_0000_0001_1111_1111_1111_1110:    data_out = 5'b1_1111; 

    default: data_out = 5'b0_0000;
    endcase
end

endmodule //decode