library verilog;
use verilog.vl_types.all;
entity tb_tdc is
end tb_tdc;
