library verilog;
use verilog.vl_types.all;
entity tb_tdc_his is
end tb_tdc_his;
